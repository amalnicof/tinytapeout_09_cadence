`timescale 1ns / 1ps

interface i2s_if;
  logic mclk;
  logic sclk;
  logic lrck;
  logic adc;
  logic dac;

  modport Slave(input mclk, input sclk, input lrck, output adc, input dac);
endinterface  // i2s_if

interface spi_if;
  logic sclk;
  logic mosi;
  logic cs;  // Active low chip-select

  modport Master(output sclk, output mosi, output cs);
endinterface

class I2SSlaveModel;
  virtual interface i2s_if.Slave i2s;

  function new(virtual interface i2s_if.Slave s);
    i2s = s;
    i2s.adc = 1'b0;
  endfunction  //new()

  task static SendAdc(input logic signed [23:0] data);
    @(posedge i2s.lrck);  // Only send data on high lrck

    for (int i = 0; i < 24; i++) begin
      @(negedge i2s.sclk);
      i2s.adc = data[23-i];
    end
  endtask

  task static ReadDac(output logic signed [23:0] data);
    @(posedge i2s.lrck);  // Only read data on high lrck
    @(posedge i2s.sclk);  // Skip first sample pulse

    for (int i = 0; i < 24; i++) begin
      @(posedge i2s.sclk);
      data = {data[22:0], i2s.dac};
    end
  endtask
endclass  // I2SSlaveModel

class SPIMasterModel;
  virtual interface spi_if.Master spi;
  logic stopClockGen;

  function new(virtual interface spi_if.Master s);
    spi = s;
    spi.sclk = 1'b0;
    spi.mosi = 1'b0;
    spi.cs = 1'b1;
  endfunction

  task static GenerateClock();
    // Generate 1MHz clock
    while (!stopClockGen) begin
      #500ns;
      spi.sclk = !spi.sclk;
    end
  endtask  // static

  task static SendData(input logic data[]);
    stopClockGen = 0;

    fork
      GenerateClock();
      begin
        @(posedge spi.sclk);
        spi.cs = 1'b0;

        for (int i = 0; i < data.size; i++) begin
          @(negedge spi.sclk);
          spi.mosi = data[i];
        end

        @(negedge spi.sclk);
        spi.cs = 1'b1;
        stopClockGen = 1'b1;
      end
    join
  endtask  // static
endclass

module tb_FIREngine ();
  localparam integer NTaps = 9;
  localparam integer NCoeff = (NTaps + 1) / 2;

  logic signed [11:0] expFilterOutput;
  logic signed [23:0] adcData;
  logic signed [23:0] dacData;

  i2s_if i2s ();
  spi_if spi ();
  I2SSlaveModel i2sModel;
  SPIMasterModel spiModel;

  // Configuration
  logic symCoeffs;
  logic [3:0] clockConfig;
  logic signed [11:0] coeffs[NCoeff];
  logic configData[1+4+(12*NCoeff)];

  // DUT signals
  logic clk;
  logic reset;

  FIREngine #(
      .NTaps(NTaps)
  ) dut (
      .clk(clk),
      .reset(reset),
      .mclk(i2s.mclk),
      .sclk(i2s.sclk),
      .lrck(i2s.lrck),
      .adc(i2s.adc),
      .dac(i2s.dac),
      .spiClk(spi.sclk),
      .mosi(spi.mosi),
      .cs(spi.cs)
  );

  task static WaitClock(input int cycles);
    repeat (cycles) @(posedge clk);
  endtask  // static

  task static ComputeFilterResponse(input logic [11:0] in, output logic [11:0] out);
    static logic signed [11:0] filterSamples[NTaps] = '{NTaps{12'd0}};
    logic signed [24:0] acc;

    logic signed [12:0] outInt;

    begin
      filterSamples = {in, filterSamples[0:NTaps-2]};
      acc = 0;
      for (int i = 0; i < NCoeff - 1; i++) begin
        if (symCoeffs) begin
          acc += (filterSamples[i] + filterSamples[NTaps-1-i]) * coeffs[i];
        end else begin
          acc += (filterSamples[i] - filterSamples[NTaps-1-i]) * coeffs[i];
        end
      end
      acc += coeffs[NCoeff-1] * filterSamples[NTaps/2];

      // Convert to output format
      outInt = acc >>> 11;
      if (outInt > signed'(13'h7ff)) begin
        out = 12'h7ff;
      end else if (outInt < signed'(12'h800)) begin
        out = signed'(12'h800);
      end else begin
        out = outInt[11:0];
      end
    end

  endtask  // static

  // Generate 32MHz clock
  initial begin
    clk = 0;
    forever begin
      #15.625 clk = ~clk;
    end
  end

  initial begin
    $dumpfile("outputs/tb_FIREngine_trace.vcd");
    $dumpvars(0, tb_FIREngine);

    $display("===================");
    $display("FIREngine Testbench");
    $display("===================");

    i2sModel = new(i2s.Slave);
    spiModel = new(spi.Master);

    // Reset core
    reset = 1;
    WaitClock(3);
    reset = 0;
    WaitClock(2);

    // Test configuration
    $display("Test configuration");
    symCoeffs   = 1'b1;
    clockConfig = $urandom();
    for (int i = 0; i < NCoeff; i++) begin
      coeffs[i] = $urandom() & 12'h7ff;
    end
    configData = {>>{{<<12{coeffs}}, symCoeffs, clockConfig}};
    spiModel.SendData(configData);

    assert (clockConfig == dut.clockConfig)
    else $error("clockConfig incorrect, should be %h not %h", clockConfig, dut.clockConfig);
    for (int i = 0; i < NCoeff; i++) begin
      assert (coeffs[i] == dut.firInst.coeffs[i])
      else
        $error("coeff incorrect, at %d should be %h not %h", i, coeffs[i], dut.firInst.coeffs[i]);
    end

    $display("Test impulse response");
    symCoeffs = 1'b1;
    clockConfig = 4'd0;
    dut.configStore.shiftReg = {symCoeffs, clockConfig};
    dut.firInst.samples = '{NTaps{12'd0}};

    adcData = 1'b1 << 22;
    i2sModel.SendAdc(adcData);
    for (int i = 0; i < NTaps + 1; i++) begin
      ComputeFilterResponse(i == 0 ? adcData >>> 12 : 0, expFilterOutput);
      i2sModel.ReadDac(dacData);

      assert (dacData == {expFilterOutput, 12'b0})
      else
        $error(
            "Impulse response incorrect, at %d should be %h not %h",
            i,
            {
              expFilterOutput, 12'b0
            },
            dacData
        );
    end

    $display("Test random data response");
    adcData = $urandom();
    i2sModel.SendAdc(adcData);
    for (int i = 0; i < NTaps * 2; i++) begin
      fork
        begin
          ComputeFilterResponse(adcData >>> 12, expFilterOutput);
          adcData = $urandom();
          i2sModel.SendAdc(adcData);
        end
        begin
          i2sModel.ReadDac(dacData);
        end
      join

      assert (dacData == {expFilterOutput, 12'b0})
      else
        $error(
            "Response incorrect, at %d should be %h not %h", i, {expFilterOutput, 12'b0}, dacData
        );
    end

    for (int i = 0; i < NTaps + 1; i++) begin
      fork
        begin
          ComputeFilterResponse(adcData >>> 12, expFilterOutput);
          adcData = 0;
          i2sModel.SendAdc(0);
        end
        begin
          i2sModel.ReadDac(dacData);
        end
      join

      assert (dacData == {expFilterOutput, 12'b0})
      else
        $error(
            "Fading response incorrect, at %d should be %h not %h",
            i,
            {
              expFilterOutput, 12'b0
            },
            dacData
        );
    end

    $display("Test anti-symmetric impulse");
    symCoeffs = 1'b0;
    dut.configStore.shiftReg = {symCoeffs, clockConfig};
    dut.firInst.samples = '{NTaps{12'd0}};

    adcData = 1'b1 << 11;
    i2sModel.SendAdc(adcData);
    for (int i = 0; i < NTaps + 1; i++) begin
      ComputeFilterResponse(i == 0 ? adcData >>> 12 : 0, expFilterOutput);
      i2sModel.ReadDac(dacData);

      assert (dacData == {expFilterOutput, 12'b0})
      else
        $error(
            "Anti-Sym, Impulse response incorrect, at %d should be %h not %h",
            i,
            {
              expFilterOutput, 12'b0
            },
            dacData
        );
    end

    WaitClock(16);
    $display("Testing complete.");
    $display("=================");
    $finish();
  end
endmodule
