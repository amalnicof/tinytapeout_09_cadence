/*
 * Module `fir`
 *
 * FIR Filter
 * Coefficients have the format SFix<1,m>, where m is DataWidth-1. For 12 bit data, the format is 1
 * sign bit and 11 fractional bits.
 * Input and output samples are unsigned integers of size DataWidth.
 */


`timescale 1ns / 1ps

module fir #(
    parameter integer DataWidth = 12,
    parameter integer NTaps = 8,

    localparam integer NCoeffs = NTaps / 2,
    localparam integer AccumulatorWidth = $clog2(
        ((1 << DataWidth) - 1) * NTaps
    ) + DataWidth - 1 + 1  // max int + frac + sign
) (
    input wire clk,
    input wire rst,
    input wire start,
    input wire lock,  // lock signal to stop coefficient shifting
    output logic done,  // Done pulse when output data is valid
    input wire coeff_load_in,
    input wire coeff_in,  // Coefficients, SFix<1,11>
    input wire [DataWidth-1:0] x,  // Input samples UFix<12,0>
    output logic [DataWidth-1:0] y  // Output samples UFix<12,0>
);
  generate
    if (NTaps % 2 == 1) begin : g_ParameterVerification_NTaps
      $fatal("NTaps must be even.");
    end
  endgenerate

  localparam integer SAMPLE_CNT_BITS = $clog2(NCoeffs);
  localparam integer BITS_CNT_BITS = $clog2(DataWidth);

  // control signals
  logic sft, sample_cnt_en, bit_cnt_en, mac_en, sample_cnt_rst;

  // samples LSFR
  // When a new sample is shifted in, the entire LSFR advances.
  // During the MAC operation, the LSFR is split in half, and advances in opposite directions.
  // This allows the MAC process to just select from the LSB and MSB of the entire lsfr
  logic [DataWidth-1:0] samples[NTaps];
  always_ff @(posedge clk) begin
    if (rst) begin
      // reset
      samples <= '{NTaps{DataWidth'(0)}};
    end else begin
      // shifting
      if (start) begin
        // Shift in new sample
        samples <= {x, samples[0:NTaps-2]};
      end else if (sft) begin
        // Split the LSFR in 2
        // x1 x2 x3 x4 | x5 x6 x7 x8
        // x2 x3 x4 x1 | x8 x5 x6 x7
        // x3 x4 x1 x2 | x7 x8 x5 x6
        // ...
        samples <= {samples[1:(NTaps/2)-1], samples[0], samples[NTaps-1], samples[NTaps/2:NTaps-2]};
      end
    end
  end

  integer k;
  integer f;
  // coefficients LSFR
  // When loading coefficients, it becomes a bit lsfr, where the new bit is shifted from the LSB
  // During the MAC operation, it shifts by DataWidth downwards
  reg [DataWidth-1:0] coeffs[NCoeffs];
  always_ff @(posedge clk) begin
    if (rst) begin
      // reset
      coeffs <= '{NCoeffs{DataWidth'(0)}};
    end else begin
      // shifting
      if (coeff_load_in) begin
        coeffs[0][0] <= coeff_in;
        for (k = 0; k < NCoeffs - 1; k++) begin
          // connection between coeffs
          coeffs[k+1][0] <= coeffs[k][DataWidth-1];

          // Connection within coeffs
          for (f = 0; f < DataWidth - 1; f++) begin
            coeffs[k][f+1] <= coeffs[k][f];
          end
        end

        // Connection within last coeff
        for (f = 0; f < DataWidth - 1; f++) begin
          coeffs[NCoeffs-1][f+1] <= coeffs[NCoeffs-1][f];
        end
      end else if (sft && !lock) begin
        coeffs <= {coeffs[1:NCoeffs-1], coeffs[0]};
      end
    end
  end

  // sample counter
  reg [SAMPLE_CNT_BITS-1:0] sample_cnt;
  always_ff @(posedge clk) begin
    if (rst) begin
      sample_cnt <= 'd0;
    end else begin
      if (sample_cnt_en) begin
        sample_cnt <= sample_cnt + 1'b1;
      end else if (sample_cnt_rst) begin
        sample_cnt <= 'd0;
      end
    end
  end

  // bit counter
  reg [BITS_CNT_BITS-1:0] bit_cnt;
  always_ff @(posedge clk) begin
    if (rst) begin
      bit_cnt <= 'd0;
    end else begin
      if ((bit_cnt_en == 1'b1) && (bit_cnt < DataWidth - 1)) begin
        bit_cnt <= bit_cnt + 1'b1;
      end else begin
        bit_cnt <= 'd0;
      end
    end
  end

  // MAC: Multiply and Accumulate
  logic [1:0] sel;
  logic [AccumulatorWidth-1:0] currCoeff;
  logic [AccumulatorWidth-1:0] currCoeff2;
  logic [AccumulatorWidth-1:0] mux_out;
  logic [AccumulatorWidth-1:0] acc_in;
  logic [AccumulatorWidth-1:0] accQ;
  always_comb begin
    // create select signal through filter symmetry
    sel = samples[0][bit_cnt] + samples[NTaps-1][bit_cnt];
    currCoeff = coeffs[0] << bit_cnt;
    currCoeff2 = currCoeff << 1;
    // MUX
    case (sel)
      2'b00:   mux_out = 'd0;
      2'b01:   mux_out = currCoeff;
      2'b10:   mux_out = currCoeff2;
      default: mux_out = 'd0;
    endcase
    acc_in = accQ + mux_out;
  end

  // accumulator register
  always_ff @(posedge clk) begin
    if (rst) begin
      accQ <= 'd0;
    end else begin
      if (start) begin
        accQ <= 'd0;
      end else if (mac_en) begin
        accQ <= acc_in;
      end
    end
  end

  // Output value
  always_comb begin
    // Convert from SFix to UFix, TODO IMP SIGN
    y = (accQ >> (DataWidth - 1)) & 12'hfff;  // Remove fractional bits, truncate to DataWidth
  end

  // STATE MACHINE
  typedef enum logic [1:0] {
    IDLE,
    COEFF_LD,
    OP,
    SHIFT
  } state_e;

  state_e n_state, state;
  // transition states
  always_ff @(posedge clk) begin
    if (rst) begin
      state <= IDLE;
    end else begin
      state <= n_state;

      if (state == SHIFT && n_state == IDLE) begin
        done <= 1'b1;
      end else begin
        done <= 1'b0;
      end
    end
  end

  // next state
  always_comb begin
    case (state)
      IDLE: begin
        if (start) n_state = OP;
        else if (coeff_load_in) n_state = COEFF_LD;
        else n_state = IDLE;
      end

      COEFF_LD: begin
        if (coeff_load_in) n_state = COEFF_LD;
        else n_state = IDLE;
      end

      OP: begin
        if (bit_cnt < DataWidth - 2) n_state = OP;
        else n_state = SHIFT;
      end

      SHIFT: begin
        if (sample_cnt < NCoeffs - 1) n_state = OP;
        else n_state = IDLE;
      end

      default: begin
      end
    endcase
  end

  // control signals
  always_comb begin
    sft = 1'b0;
    sample_cnt_en = 1'b0;
    bit_cnt_en = 1'b0;
    mac_en = 1'b0;
    sample_cnt_rst = 1'b0;
    case (state)
      IDLE: begin
        sample_cnt_rst = 1'b1;
      end

      COEFF_LD: begin
      end

      OP: begin
        mac_en = 1'b1;
        bit_cnt_en = 1'b1;
      end

      SHIFT: begin
        sft = 1'b1;
        mac_en = 1'b1;
        bit_cnt_en = 1'b1;
        sample_cnt_en = 1'b1;
      end

      default: begin
      end
    endcase
  end
endmodule
